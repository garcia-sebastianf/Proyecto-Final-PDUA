LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------
ENTITY uProgramMemory IS
PORT(	uaddr	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
		UI		: 	OUT 	STD_LOGIC_VECTOR(28 DOWNTO 0));
END ENTITY uProgramMemory;
-----------------------------------------------------
ARCHITECTURE behavioral OF uProgramMemory IS
BEGIN
	
	MUI: PROCESS(uaddr)
	BEGIN
		CASE uaddr IS
	-- Complete the following values according to your particular implementation 
	-- Unused postions do not affect the operation of the ROM
			-- FETCH 							    
			WHEN "00000000" => UI <= "00000000000001000001110001001"; 
			WHEN "00000001" => UI <= "01100000000010000001110000000"; 
			WHEN "00000010" => UI <= "00000000000000100001110000000"; 
			WHEN "00000011" => UI <= "00000000000000010001010001000"; 
																					
			--00001	 MOV ACC,A 
			WHEN "00001000" => UI <= "10000001111110000001110001000";

			--00010  MOV A,ACC
			WHEN "00010000" => UI <= "10000011101110000001110001000";

			--00011	 MOV ACC,CTE 
			WHEN "00011000" => UI <= "00000000000001000000010000000";
			WHEN "00011001" => UI <= "01100000000010000000010000000";
			WHEN "00011010" => UI <= "00000000000000100000010000000";
			WHEN "00011011" => UI <= "00000000011110010001110001000";

			--00100  MOV ACC,[DPTR]
			WHEN "00100000" => UI <= "00000001000001000000010000000";
			WHEN "00100001" => UI <= "00000000000000000000010000000";
			WHEN "00100010" => UI <= "00000000000000100000010000000";
			WHEN "00100011" => UI <= "00000000011110010001110001000";

			--00101  MOV DPTR,ACC
			WHEN "00101000" => UI <= "10000011101010000001110001000";
		
			-- 00110 MOV [DPTR],ACC	
			WHEN "00110000" => UI <= "00000001000001000000010000000";
			WHEN "00110001" => UI <= "10000011100000100000010000000";
         WHEN "00110010" => UI <= "00000000000000000011110001000";

			 -- 01000 AND ACC,A	 
			WHEN "01000000" => UI <= "10100001111110000001110001000";

			 -- 10000 OR ACC,A	
			WHEN "10000000" => UI <= "10110001111110000001110001000";
			
			 -- 10001 XOR ACC,A	
			WHEN "10001000" => UI <= "11000001111110000001110001000";

			-- 01001 ADD ACC,A
			WHEN "01001000" => UI <= "11010001111110000001110001000";

			-- 10010 INC ACC
			WHEN "10010000" => UI <= "11100011111110000001110001000";

			-- 00111 INV ACC
			WHEN "00111000" => UI <= "10010011111110000001110001000";
			
			-- 00111 NEG ACC
			WHEN "10011000" => UI <= "11110011111110000001110001000";

			-- 10100 SLL ACC
			WHEN "10100000" => UI <= "10001011111110000001110001000";
			
			-- 10101 SLR ACC
			WHEN "10101000" => UI <= "10000111111110000001110001000";			
			
			-- 01010 JMP CTE
			WHEN "01010000" => UI <= "00000000000001000000010000000";
			WHEN "01010001" => UI <= "01100000000010000000010000000";
			WHEN "01010010" => UI <= "00000000000000100000010000000";
			WHEN "01010011" => UI <= "00000000000010010001110001000";
			
			-- 01011 JZ 
			WHEN "01011000" => UI <= "00000000000000000000010010010";
			WHEN "01011001" => UI <= "01100000000010000001110001000";
			WHEN "01011010" => UI <= "00000000000001000000010000000";
			WHEN "01011011" => UI <= "01100000000010000000010000000";
			WHEN "01011100" => UI <= "00000000000000100000010000000";
			WHEN "01011101" => UI <= "00000000000010010001110001000";

			-- 01100 JN 
			WHEN "01100000" => UI <= "00000000000000000000010011010";
			WHEN "01100001" => UI <= "01100000000010000001110001000";
			WHEN "01100010" => UI <= "00000000000001000000010000000";
			WHEN "01100011" => UI <= "01100000000010000000010000000";
			WHEN "01100100" => UI <= "00000000000000100000010000000";
			WHEN "01100101" => UI <= "00000000000010010001110001000";
			
			-- 01101 JC 
			WHEN "01101000" => UI <= "00000000000000000000010100010";
			WHEN "01101001" => UI <= "01100000000010000001110001000";
			WHEN "01101010" => UI <= "00000000000001000000010000000";
			WHEN "01101011" => UI <= "01100000000010000000010000000";
			WHEN "01101100" => UI <= "00000000000000100000010000000";
			WHEN "01101101" => UI <= "00000000000010010001110001000";
			
			--11111 HALT 
			WHEN "11111000" => UI <= "00000000000000000000011000000";
			
			WHEN others => UI <= (others => 'X');
		END CASE;
	END PROCESS;
END ARCHITECTURE Behavioral;